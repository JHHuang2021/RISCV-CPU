module Fetcher(
    input wire clk,
    input wire rst,
    input wire rdy,

);

endmodule